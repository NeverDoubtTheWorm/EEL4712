library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity alu_ns_tb is
end alu_ns_tb;

architecture TB of alu_ns_tb is

  component alu_ns

    generic (
      WIDTH    :     positive := 16
      );
    port (
      input1   : in  std_logic_vector(WIDTH-1 downto 0);
      input2   : in  std_logic_vector(WIDTH-1 downto 0);
      sel      : in  std_logic_vector(3 downto 0);
      output   : out std_logic_vector(WIDTH-1 downto 0);
      overflow : out std_logic
      );

  end component;

  constant WIDTH    : positive                           := 8;
  signal   input1   : std_logic_vector(WIDTH-1 downto 0) := (others => '0');
  signal   input2   : std_logic_vector(WIDTH-1 downto 0) := (others => '0');
  signal   sel      : std_logic_vector(3 downto 0)       := (others => '0');
  signal   output   : std_logic_vector(WIDTH-1 downto 0);
  signal   overflow : std_logic;

begin  -- TB

  UUT : alu_ns
    generic map (WIDTH => WIDTH)
    port map (
      input1           => input1,
      input2           => input2,
      sel              => sel,
      output           => output,
      overflow         => overflow);


  process

    function sum_test (
      constant input1      : integer;
      constant input2      : integer)
      return std_logic_vector is
    begin
      return std_logic_vector(to_unsigned((input1+input2) mod 65536, WIDTH));
    end sum_test;
	 
    function sub_test (
      constant input1      : integer;
      constant input2      : integer)
      return std_logic_vector is
    begin
      return std_logic_vector(to_unsigned((input1-input2) mod 65536, WIDTH));
    end sub_test;

    function MULOFL_test (
      constant input1      : integer;
      constant input2      : integer;
      constant select	   : integer)
      return std_logic is
    begin
      if (input1*input2 > "11111111") then
        return '1';
      else
        return '0';
      end if;
    end carry_test;
	 
  begin

    -- test 2+6 (no overflow)
    sel    <= "0000";
    input1 <= conv_std_logic_vector(2, input1'length);
    input2 <= conv_std_logic_vector(6, input2'length);
    wait for 40 ns;
    assert(output = conv_std_logic_vector(8, output'length)) report "Error : 2+6 = " & integer'image(conv_integer(output)) & " instead of 8" severity warning;
    assert(overflow = '0') report "Error                                   : overflow incorrect for 2+8" severity warning;

    -- test 250+50 (with overflow)
    sel    <= "0000";
    input1 <= conv_std_logic_vector(250, input1'length);
    input2 <= conv_std_logic_vector(50, input2'length);
    wait for 40 ns;
    assert(output = conv_std_logic_vector(300, output'length)) report "Error : 250+50 = " & integer'image(conv_integer(output)) & " instead of 44" severity warning;
    assert(overflow = '1') report "Error                                     : overflow incorrect for 250+50" severity warning;

    -- test 5*6
    sel    <= "0010";
    input1 <= conv_std_logic_vector(5, input1'length);
    input2 <= conv_std_logic_vector(6, input2'length);
    wait for 40 ns;
    assert(output = conv_std_logic_vector(30, output'length)) report "Error : 5*6 = " & integer'image(conv_integer(output)) & " instead of 30" severity warning;
    assert(overflow = '0') report "Error                                    : overflow incorrect for 5*6" severity warning;

    -- test 50*60
    sel    <= "0010";
    input1 <= conv_std_logic_vector(64, input1'length);
    input2 <= conv_std_logic_vector(64, input2'length);
    wait for 40 ns;
    assert(output = conv_std_logic_vector(4096, output'length)) report "Error : 64*64 = " & integer'image(conv_integer(output)) & " instead of 0" severity warning;
    assert(overflow = '1') report "Error                                      : overflow incorrect for 64*64" severity warning;

    -- add many more tests

    wait;

  end process;



end TB;
