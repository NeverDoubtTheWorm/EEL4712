library ieee;
use ieee.std_logic_1164.all;

package lib is

-----------------------------------------------------------------------------
-- reg_en
constant accu_reg_en: std_logic_vector := "10000000000";
constant ir_reg_en	: std_logic_vector := "01000000000";
constant data_reg_en: std_logic_vector := "00100000000";
constant xh_reg_en	: std_logic_vector := "00010000000";
constant xl_reg_en	: std_logic_vector := "00001000000";
constant pch_reg_en	: std_logic_vector := "00000100000";
constant pcl_reg_en	: std_logic_vector := "00000010000";
constant arh_reg_en	: std_logic_vector := "00000001000";
constant arl_reg_en	: std_logic_vector := "00000000100";
constant sph_reg_en	: std_logic_vector := "00000000010";
constant spl_reg_en	: std_logic_vector := "00000000001";
constant none		: std_Logic_vector := "00000000000";		
-----------------------------------------------------------------------------
--Status reg en
constant carry		: std_logic_vector := "1000";
constant overflow	: std_logic_vector := "0100";
constant sign		: std_logic_vector := "0010";
constant zero		: std_logic_vector := "0001";
constant none1		: std_logic_vector := "0000";
-----------------------------------------------------------------------------
--Internal BUS sel
constant outALU		: std_logic_vector	:= "0001";
constant outACCU	: std_logic_vector 	:= "0010";
constant outDATA	: std_logic_vector 	:= "0011";
constant outXh		: std_logic_vector 	:= "0100";
constant outXl		: std_logic_vector 	:= "0101";
constant outSPh		: std_logic_vector 	:= "0110";
constant outSPl		: std_logic_vector 	:= "0111";
constant outPCh		: std_logic_vector 	:= "1000";
constant outPCl		: std_logic_vector 	:= "1001";
constant databusin	: std_logic_vector	:= "1010";
constant outIR		: std_logic_Vector 	:= "1011";
constant outAR 		: std_logic_vector	:= "1100";
-----------------------------------------------------------------------------
--BUS sel
constant internal	: std_logic_vector	:= "0001";
constant ram		: std_logic_vector 	:= "0010";
constant dip		: std_logic_vector 	:= "0011";
constant dip2		: std_logic_vector 	:= "0100";
-----------------------------------------------------------------------------
--PC ADD
constant zero2	: std_logic_vector := "000";
constant one	: std_logic_vector := "001";
constant two	: std_logic_vector := "010";	
constant three	: std_logic_vector := "011";
constant minus	: std_logic_vector := "100";
end lib;